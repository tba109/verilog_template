///////////////////////////////////////////////////////////////////////////////////////////////////////////////////
// <NAME> <DATE>
//
// <MODULE NAME>.v
//
// <DESCRIPTION> 
//////////////////////////////////////////////////////////////////////////////////////////////////////////////////

`timescale 1ns/1ns

///////////////////////////////////////////////////////////////////////////////////////////////////
// Test cases
///////////////////////////////////////////////////////////////////////////////////////////////////
`define <TEST_CASE_NAME>

module <MODULE_NAME_TB>;
   
   //////////////////////////////////////////////////////////////////////
   // I/O
   //////////////////////////////////////////////////////////////////////   
   parameter SYSCLK_PERIOD = <PERIOD_NS>;
   reg SYSCLK;
   reg SYSRESET;

   // Connections
   wire w1; 
   reg 	r1; 

   //////////////////////////////////////////////////////////////////////
   // Clock Driver
   //////////////////////////////////////////////////////////////////////
   always @(SYSCLK)
     #(SYSCLK_PERIOD / 2.0) SYSCLK <= !SYSCLK;
				   
   //////////////////////////////////////////////////////////////////////
   // Simulated interfaces
   //////////////////////////////////////////////////////////////////////   
      
   //////////////////////////////////////////////////////////////////////
   // UUT
   //////////////////////////////////////////////////////////////////////   
      
   //////////////////////////////////////////////////////////////////////
   // Testbench
   //////////////////////////////////////////////////////////////////////   
   initial
     begin
	// Initializations
	SYSCLK = 1'b0;
	SYSRESET = 1'b1;
     end

   //////////////////////////////////////////////////////////////////////
   // Test case
   //////////////////////////////////////////////////////////////////////   
   `ifdef <TEST_CASE_NAME>
   initial
     begin
	// Reset	
	#(10 * SYSCLK_PERIOD);
	SYSRESET = 1'b0;
	#(20* SYSCLK_PERIOD);
	#(10 * DCLK_PERIOD);
	DRESET = 1'b0;
	#(20* DCLK_PERIOD);

	// Logging
	$display("");
	$display("------------------------------------------------------");
	$display("Test Case: <TEST_CASE_NAME>");

	// Stimulate UUT
     end
   `endif

   //////////////////////////////////////////////////////////////////////
   // Tasks (e.g., writing data, etc.)
   //////////////////////////////////////////////////////////////////////   
   
   
   
endmodule

// Local Variables:
// verilog-library-flags:("-y ../hdl/")
// End:
   
